package top_regs_Consts;
  localparam TOP_SIZE = 40;
  localparam ADDR_TOP_UART = 'h10;
  localparam ADDR_MASK_TOP_UART = 'h38;
  localparam TOP_UART_SIZE = 8;
  localparam ADDR_TOP_VIDEO = 'h20;
  localparam ADDR_MASK_TOP_VIDEO = 'h38;
  localparam TOP_VIDEO_SIZE = 8;
endpackage
