package video_Consts;
  localparam VIDEO_SIZE = 8;
  localparam ADDR_VIDEO_CTRL = 'h0;
  localparam VIDEO_CTRL_FB_EN_OFFSET = 0;
  localparam VIDEO_CTRL_FB_EN = 32'h1;
  localparam ADDR_VIDEO_BG_COLOR = 'h4;
  localparam VIDEO_BG_COLOR_COLOR_OFFSET = 0;
  localparam VIDEO_BG_COLOR_COLOR = 32'hffffff;
endpackage
