`default_nettype none

module Text_Generator(
    clk_i,
    rst_i,

    end_of_frame_i,
    end_of_line_i,
    hsync_n_i,
    vsync_n_i,
    visible_i,

    bg_rgb_i,
    fg_rgb_i,

    end_of_frame_o,
    end_of_line_o,
    hsync_n_o,
    vsync_n_o,
    visible_o,
    rgb_o,

    // Memory interface
    addr_o,         // address in 16-bit words
    rd_strobe_o,    // read strobe: we expect the data exactly 3 cycles after signalling this

    data_i
);

input clk_i, rst_i;
input end_of_frame_i, end_of_line_i, hsync_n_i, vsync_n_i, visible_i;
input[23:0] bg_rgb_i, fg_rgb_i;
output reg end_of_frame_o, end_of_line_o, hsync_n_o, vsync_n_o, visible_o;
output reg[23:0] rgb_o;

// 60x21 = 1260 = 11 bits
output reg[10:0] addr_o;
output reg rd_strobe_o;
input[15:0] data_i;

localparam CHAR_W = 6;
localparam CHAR_H = 11;
wire[CHAR_W-1:0] fontdata[0:96 * 11 - 1];   // FIXME: this does NOT infer a ROM!

reg[6:0] col;   // 0 to 360/6
reg[7:0] row;   // 0 to 240/11
reg[$clog2(6)-1:0] xx;
reg[$clog2(11)-1:0] yy;
reg[CHAR_W-1:0] buffer;

reg[$clog2(96 * CHAR_H - 1)-1:0] addr;
reg[$clog2(360)-1:0] x;
reg[$clog2(240)-1:0] y;

reg[6:0] char_data;

reg start_of_line;  // end_of_line_i delayed by 1 clock

always @ (posedge clk_i) begin
    if (rst_i) begin
        col <= 0;
        row <= 0;
        xx <= 0;
        yy <= 0;
        x <= 0;
        y <= 0;
    end else begin
        if (end_of_frame_i) begin
            row <= 0;
            yy <= 0;
            y <= 0;

            // TODO: how do we trigger fetch of the first character?
        end else if (end_of_line_i) begin
            if (yy < CHAR_H - 1) begin
                yy <= yy + 1;
            end else begin
                yy <= 0;
                row <= row + 1;
            end

            y <= y + 1;
        end

        addr <= char_data * 11 + yy;

        if (end_of_line_i) begin
            col <= 0;
            xx <= 0;
            x <= 0;
        end else if (visible_i) begin
            if (xx < CHAR_W - 1) begin
                xx <= xx + 1;
            end else begin
                xx <= 0;
                col <= col + 1;
            end

            buffer <= {buffer[CHAR_W-2:0], 1'b0};
            x <= x + 1;
        end

        // this needs to be done:
        //  - exactly at xx == CHAR_W-1
        //  - sometime after start_of_line and before xx = 0 && visible_i = 1
        if ((xx == 0 && !visible_i) || xx == CHAR_W - 1) begin
            buffer <= fontdata[addr];
        end
    end

    start_of_line <= end_of_line_i;

    end_of_frame_o <= end_of_frame_i;
    end_of_line_o <= end_of_line_i;
    hsync_n_o <= hsync_n_i;
    vsync_n_o <= vsync_n_i;
    visible_o <= visible_i;
    rgb_o = (buffer[CHAR_W-1] ? fg_rgb_i : bg_rgb_i);
end

// Memory access control:
// We are using the "slave timing" mode of BT656_Encoder, which means we must present our data just after seeing the pre_accept strobe
// After seeing accept_o, we can start loading the next character (we wait 1 cycle to see the updated row & col)
// BT656 is 2pixels / 4clk at 27 MHz. With 6-pixel characters, we get 12 clk per char
localparam MEM_IDLE = 0;
localparam MEM_STROBE_RD = 1;
localparam MEM_DATA_READY = 4;

reg[2:0] mem_state;

always @ (posedge clk_i) begin
    rd_strobe_o <= 1'b0;

    if (rst_i) begin
        mem_state <= MEM_IDLE;
        addr_o <= 0;
        char_data <= 0;
    end else begin
        // $display("begin cycle: x=%d, yy=%d, acc=%d, p_a=%d, sol=%d", x, yy, accept_i, pre_accept_i, start_of_line_i);

        if (start_of_line) begin
            addr_o <= row * 60;
            char_data <= row * 1;
        end

        // if (accept_i && xx == 0) begin
        //     $display("state=%d at 1st acc (x=%d, xx=0)", mem_state, x);
        // end

        if (mem_state == MEM_IDLE) begin
            if ((visible_i && xx == 0) || start_of_line) begin
                // $display("MEM_IDLE: begin read cycle at r,c %d,%d; acc=%d, sol=%d", row, col, accept_i, start_of_line_i);
                mem_state <= MEM_STROBE_RD;
            end

            if (visible_i && xx == 0) begin
                addr_o <= addr_o + 1;
                char_data <= char_data + 1;
                // $display("inc char_data to %d at x=%d", char_data + 1, x);
            end
        end else if (mem_state == MEM_STROBE_RD) begin
            // $display("MEM_STROBE_RD: read addr %d while row=%d, col=%d, x=%d", addr_o, row, col, x);
            rd_strobe_o <= 1'b1;
        end else if (mem_state == MEM_DATA_READY) begin
            // char_data <= data_i;
        end

        if (mem_state == MEM_DATA_READY) begin
            // $display("x=%d, mem_state=%d", x, mem_state);
            mem_state <= 0;
        end else if (mem_state > 0) begin
            // $display("x=%d, mem_state=%d", x, mem_state);
            mem_state <= mem_state + 1'b1;
        end
    end
end

assign fontdata[ 0 * 11 +  0] = 6'b000000;
assign fontdata[ 0 * 11 +  1] = 6'b000000;
assign fontdata[ 0 * 11 +  2] = 6'b000000;
assign fontdata[ 0 * 11 +  3] = 6'b000000;
assign fontdata[ 0 * 11 +  4] = 6'b000000;
assign fontdata[ 0 * 11 +  5] = 6'b000000;
assign fontdata[ 0 * 11 +  6] = 6'b000000;
assign fontdata[ 0 * 11 +  7] = 6'b000000;
assign fontdata[ 0 * 11 +  8] = 6'b000000;
assign fontdata[ 0 * 11 +  9] = 6'b000000;
assign fontdata[ 0 * 11 + 10] = 6'b000000;
assign fontdata[ 1 * 11 +  0] = 6'b000000;
assign fontdata[ 1 * 11 +  1] = 6'b001000;
assign fontdata[ 1 * 11 +  2] = 6'b001000;
assign fontdata[ 1 * 11 +  3] = 6'b001000;
assign fontdata[ 1 * 11 +  4] = 6'b001000;
assign fontdata[ 1 * 11 +  5] = 6'b001000;
assign fontdata[ 1 * 11 +  6] = 6'b001000;
assign fontdata[ 1 * 11 +  7] = 6'b000000;
assign fontdata[ 1 * 11 +  8] = 6'b001000;
assign fontdata[ 1 * 11 +  9] = 6'b000000;
assign fontdata[ 1 * 11 + 10] = 6'b000000;
assign fontdata[ 2 * 11 +  0] = 6'b000000;
assign fontdata[ 2 * 11 +  1] = 6'b010100;
assign fontdata[ 2 * 11 +  2] = 6'b010100;
assign fontdata[ 2 * 11 +  3] = 6'b010100;
assign fontdata[ 2 * 11 +  4] = 6'b000000;
assign fontdata[ 2 * 11 +  5] = 6'b000000;
assign fontdata[ 2 * 11 +  6] = 6'b000000;
assign fontdata[ 2 * 11 +  7] = 6'b000000;
assign fontdata[ 2 * 11 +  8] = 6'b000000;
assign fontdata[ 2 * 11 +  9] = 6'b000000;
assign fontdata[ 2 * 11 + 10] = 6'b000000;
assign fontdata[ 3 * 11 +  0] = 6'b000000;
assign fontdata[ 3 * 11 +  1] = 6'b010100;
assign fontdata[ 3 * 11 +  2] = 6'b010100;
assign fontdata[ 3 * 11 +  3] = 6'b111110;
assign fontdata[ 3 * 11 +  4] = 6'b010100;
assign fontdata[ 3 * 11 +  5] = 6'b111110;
assign fontdata[ 3 * 11 +  6] = 6'b010100;
assign fontdata[ 3 * 11 +  7] = 6'b010100;
assign fontdata[ 3 * 11 +  8] = 6'b000000;
assign fontdata[ 3 * 11 +  9] = 6'b000000;
assign fontdata[ 3 * 11 + 10] = 6'b000000;
assign fontdata[ 4 * 11 +  0] = 6'b000000;
assign fontdata[ 4 * 11 +  1] = 6'b001000;
assign fontdata[ 4 * 11 +  2] = 6'b011100;
assign fontdata[ 4 * 11 +  3] = 6'b101010;
assign fontdata[ 4 * 11 +  4] = 6'b101000;
assign fontdata[ 4 * 11 +  5] = 6'b011100;
assign fontdata[ 4 * 11 +  6] = 6'b001010;
assign fontdata[ 4 * 11 +  7] = 6'b101010;
assign fontdata[ 4 * 11 +  8] = 6'b011100;
assign fontdata[ 4 * 11 +  9] = 6'b001000;
assign fontdata[ 4 * 11 + 10] = 6'b000000;
assign fontdata[ 5 * 11 +  0] = 6'b000000;
assign fontdata[ 5 * 11 +  1] = 6'b000000;
assign fontdata[ 5 * 11 +  2] = 6'b010010;
assign fontdata[ 5 * 11 +  3] = 6'b101010;
assign fontdata[ 5 * 11 +  4] = 6'b010100;
assign fontdata[ 5 * 11 +  5] = 6'b001000;
assign fontdata[ 5 * 11 +  6] = 6'b010100;
assign fontdata[ 5 * 11 +  7] = 6'b101010;
assign fontdata[ 5 * 11 +  8] = 6'b100100;
assign fontdata[ 5 * 11 +  9] = 6'b000000;
assign fontdata[ 5 * 11 + 10] = 6'b000000;
assign fontdata[ 6 * 11 +  0] = 6'b000000;
assign fontdata[ 6 * 11 +  1] = 6'b000000;
assign fontdata[ 6 * 11 +  2] = 6'b011000;
assign fontdata[ 6 * 11 +  3] = 6'b100100;
assign fontdata[ 6 * 11 +  4] = 6'b101000;
assign fontdata[ 6 * 11 +  5] = 6'b010000;
assign fontdata[ 6 * 11 +  6] = 6'b101010;
assign fontdata[ 6 * 11 +  7] = 6'b100100;
assign fontdata[ 6 * 11 +  8] = 6'b011010;
assign fontdata[ 6 * 11 +  9] = 6'b000000;
assign fontdata[ 6 * 11 + 10] = 6'b000000;
assign fontdata[ 7 * 11 +  0] = 6'b000000;
assign fontdata[ 7 * 11 +  1] = 6'b001000;
assign fontdata[ 7 * 11 +  2] = 6'b001000;
assign fontdata[ 7 * 11 +  3] = 6'b001000;
assign fontdata[ 7 * 11 +  4] = 6'b000000;
assign fontdata[ 7 * 11 +  5] = 6'b000000;
assign fontdata[ 7 * 11 +  6] = 6'b000000;
assign fontdata[ 7 * 11 +  7] = 6'b000000;
assign fontdata[ 7 * 11 +  8] = 6'b000000;
assign fontdata[ 7 * 11 +  9] = 6'b000000;
assign fontdata[ 7 * 11 + 10] = 6'b000000;
assign fontdata[ 8 * 11 +  0] = 6'b000000;
assign fontdata[ 8 * 11 +  1] = 6'b000100;
assign fontdata[ 8 * 11 +  2] = 6'b001000;
assign fontdata[ 8 * 11 +  3] = 6'b001000;
assign fontdata[ 8 * 11 +  4] = 6'b010000;
assign fontdata[ 8 * 11 +  5] = 6'b010000;
assign fontdata[ 8 * 11 +  6] = 6'b010000;
assign fontdata[ 8 * 11 +  7] = 6'b001000;
assign fontdata[ 8 * 11 +  8] = 6'b001000;
assign fontdata[ 8 * 11 +  9] = 6'b000100;
assign fontdata[ 8 * 11 + 10] = 6'b000000;
assign fontdata[ 9 * 11 +  0] = 6'b000000;
assign fontdata[ 9 * 11 +  1] = 6'b010000;
assign fontdata[ 9 * 11 +  2] = 6'b001000;
assign fontdata[ 9 * 11 +  3] = 6'b001000;
assign fontdata[ 9 * 11 +  4] = 6'b000100;
assign fontdata[ 9 * 11 +  5] = 6'b000100;
assign fontdata[ 9 * 11 +  6] = 6'b000100;
assign fontdata[ 9 * 11 +  7] = 6'b001000;
assign fontdata[ 9 * 11 +  8] = 6'b001000;
assign fontdata[ 9 * 11 +  9] = 6'b010000;
assign fontdata[ 9 * 11 + 10] = 6'b000000;
assign fontdata[10 * 11 +  0] = 6'b000000;
assign fontdata[10 * 11 +  1] = 6'b000000;
assign fontdata[10 * 11 +  2] = 6'b000000;
assign fontdata[10 * 11 +  3] = 6'b001000;
assign fontdata[10 * 11 +  4] = 6'b101010;
assign fontdata[10 * 11 +  5] = 6'b011100;
assign fontdata[10 * 11 +  6] = 6'b101010;
assign fontdata[10 * 11 +  7] = 6'b001000;
assign fontdata[10 * 11 +  8] = 6'b000000;
assign fontdata[10 * 11 +  9] = 6'b000000;
assign fontdata[10 * 11 + 10] = 6'b000000;
assign fontdata[11 * 11 +  0] = 6'b000000;
assign fontdata[11 * 11 +  1] = 6'b000000;
assign fontdata[11 * 11 +  2] = 6'b000000;
assign fontdata[11 * 11 +  3] = 6'b001000;
assign fontdata[11 * 11 +  4] = 6'b001000;
assign fontdata[11 * 11 +  5] = 6'b111110;
assign fontdata[11 * 11 +  6] = 6'b001000;
assign fontdata[11 * 11 +  7] = 6'b001000;
assign fontdata[11 * 11 +  8] = 6'b000000;
assign fontdata[11 * 11 +  9] = 6'b000000;
assign fontdata[11 * 11 + 10] = 6'b000000;
assign fontdata[12 * 11 +  0] = 6'b000000;
assign fontdata[12 * 11 +  1] = 6'b000000;
assign fontdata[12 * 11 +  2] = 6'b000000;
assign fontdata[12 * 11 +  3] = 6'b000000;
assign fontdata[12 * 11 +  4] = 6'b000000;
assign fontdata[12 * 11 +  5] = 6'b000000;
assign fontdata[12 * 11 +  6] = 6'b000000;
assign fontdata[12 * 11 +  7] = 6'b011000;
assign fontdata[12 * 11 +  8] = 6'b011000;
assign fontdata[12 * 11 +  9] = 6'b001000;
assign fontdata[12 * 11 + 10] = 6'b010000;
assign fontdata[13 * 11 +  0] = 6'b000000;
assign fontdata[13 * 11 +  1] = 6'b000000;
assign fontdata[13 * 11 +  2] = 6'b000000;
assign fontdata[13 * 11 +  3] = 6'b000000;
assign fontdata[13 * 11 +  4] = 6'b000000;
assign fontdata[13 * 11 +  5] = 6'b111110;
assign fontdata[13 * 11 +  6] = 6'b000000;
assign fontdata[13 * 11 +  7] = 6'b000000;
assign fontdata[13 * 11 +  8] = 6'b000000;
assign fontdata[13 * 11 +  9] = 6'b000000;
assign fontdata[13 * 11 + 10] = 6'b000000;
assign fontdata[14 * 11 +  0] = 6'b000000;
assign fontdata[14 * 11 +  1] = 6'b000000;
assign fontdata[14 * 11 +  2] = 6'b000000;
assign fontdata[14 * 11 +  3] = 6'b000000;
assign fontdata[14 * 11 +  4] = 6'b000000;
assign fontdata[14 * 11 +  5] = 6'b000000;
assign fontdata[14 * 11 +  6] = 6'b000000;
assign fontdata[14 * 11 +  7] = 6'b011000;
assign fontdata[14 * 11 +  8] = 6'b011000;
assign fontdata[14 * 11 +  9] = 6'b000000;
assign fontdata[14 * 11 + 10] = 6'b000000;
assign fontdata[15 * 11 +  0] = 6'b000000;
assign fontdata[15 * 11 +  1] = 6'b000010;
assign fontdata[15 * 11 +  2] = 6'b000010;
assign fontdata[15 * 11 +  3] = 6'b000100;
assign fontdata[15 * 11 +  4] = 6'b000100;
assign fontdata[15 * 11 +  5] = 6'b001000;
assign fontdata[15 * 11 +  6] = 6'b001000;
assign fontdata[15 * 11 +  7] = 6'b010000;
assign fontdata[15 * 11 +  8] = 6'b010000;
assign fontdata[15 * 11 +  9] = 6'b100000;
assign fontdata[15 * 11 + 10] = 6'b100000;
assign fontdata[16 * 11 +  0] = 6'b000000;
assign fontdata[16 * 11 +  1] = 6'b000000;
assign fontdata[16 * 11 +  2] = 6'b011100;
assign fontdata[16 * 11 +  3] = 6'b100010;
assign fontdata[16 * 11 +  4] = 6'b100110;
assign fontdata[16 * 11 +  5] = 6'b101010;
assign fontdata[16 * 11 +  6] = 6'b110010;
assign fontdata[16 * 11 +  7] = 6'b100010;
assign fontdata[16 * 11 +  8] = 6'b011100;
assign fontdata[16 * 11 +  9] = 6'b000000;
assign fontdata[16 * 11 + 10] = 6'b000000;
assign fontdata[17 * 11 +  0] = 6'b000000;
assign fontdata[17 * 11 +  1] = 6'b000000;
assign fontdata[17 * 11 +  2] = 6'b001000;
assign fontdata[17 * 11 +  3] = 6'b011000;
assign fontdata[17 * 11 +  4] = 6'b101000;
assign fontdata[17 * 11 +  5] = 6'b001000;
assign fontdata[17 * 11 +  6] = 6'b001000;
assign fontdata[17 * 11 +  7] = 6'b001000;
assign fontdata[17 * 11 +  8] = 6'b001000;
assign fontdata[17 * 11 +  9] = 6'b000000;
assign fontdata[17 * 11 + 10] = 6'b000000;
assign fontdata[18 * 11 +  0] = 6'b000000;
assign fontdata[18 * 11 +  1] = 6'b000000;
assign fontdata[18 * 11 +  2] = 6'b011100;
assign fontdata[18 * 11 +  3] = 6'b100010;
assign fontdata[18 * 11 +  4] = 6'b000010;
assign fontdata[18 * 11 +  5] = 6'b000100;
assign fontdata[18 * 11 +  6] = 6'b001000;
assign fontdata[18 * 11 +  7] = 6'b010000;
assign fontdata[18 * 11 +  8] = 6'b111110;
assign fontdata[18 * 11 +  9] = 6'b000000;
assign fontdata[18 * 11 + 10] = 6'b000000;
assign fontdata[19 * 11 +  0] = 6'b000000;
assign fontdata[19 * 11 +  1] = 6'b000000;
assign fontdata[19 * 11 +  2] = 6'b011100;
assign fontdata[19 * 11 +  3] = 6'b100010;
assign fontdata[19 * 11 +  4] = 6'b000010;
assign fontdata[19 * 11 +  5] = 6'b001100;
assign fontdata[19 * 11 +  6] = 6'b000010;
assign fontdata[19 * 11 +  7] = 6'b100010;
assign fontdata[19 * 11 +  8] = 6'b011100;
assign fontdata[19 * 11 +  9] = 6'b000000;
assign fontdata[19 * 11 + 10] = 6'b000000;
assign fontdata[20 * 11 +  0] = 6'b000000;
assign fontdata[20 * 11 +  1] = 6'b000000;
assign fontdata[20 * 11 +  2] = 6'b000100;
assign fontdata[20 * 11 +  3] = 6'b001100;
assign fontdata[20 * 11 +  4] = 6'b010100;
assign fontdata[20 * 11 +  5] = 6'b100100;
assign fontdata[20 * 11 +  6] = 6'b111110;
assign fontdata[20 * 11 +  7] = 6'b000100;
assign fontdata[20 * 11 +  8] = 6'b000100;
assign fontdata[20 * 11 +  9] = 6'b000000;
assign fontdata[20 * 11 + 10] = 6'b000000;
assign fontdata[21 * 11 +  0] = 6'b000000;
assign fontdata[21 * 11 +  1] = 6'b000000;
assign fontdata[21 * 11 +  2] = 6'b111110;
assign fontdata[21 * 11 +  3] = 6'b100000;
assign fontdata[21 * 11 +  4] = 6'b111100;
assign fontdata[21 * 11 +  5] = 6'b000010;
assign fontdata[21 * 11 +  6] = 6'b000010;
assign fontdata[21 * 11 +  7] = 6'b100010;
assign fontdata[21 * 11 +  8] = 6'b011100;
assign fontdata[21 * 11 +  9] = 6'b000000;
assign fontdata[21 * 11 + 10] = 6'b000000;
assign fontdata[22 * 11 +  0] = 6'b000000;
assign fontdata[22 * 11 +  1] = 6'b000000;
assign fontdata[22 * 11 +  2] = 6'b011100;
assign fontdata[22 * 11 +  3] = 6'b100000;
assign fontdata[22 * 11 +  4] = 6'b111100;
assign fontdata[22 * 11 +  5] = 6'b100010;
assign fontdata[22 * 11 +  6] = 6'b100010;
assign fontdata[22 * 11 +  7] = 6'b100010;
assign fontdata[22 * 11 +  8] = 6'b011100;
assign fontdata[22 * 11 +  9] = 6'b000000;
assign fontdata[22 * 11 + 10] = 6'b000000;
assign fontdata[23 * 11 +  0] = 6'b000000;
assign fontdata[23 * 11 +  1] = 6'b000000;
assign fontdata[23 * 11 +  2] = 6'b111110;
assign fontdata[23 * 11 +  3] = 6'b000010;
assign fontdata[23 * 11 +  4] = 6'b000100;
assign fontdata[23 * 11 +  5] = 6'b000100;
assign fontdata[23 * 11 +  6] = 6'b001000;
assign fontdata[23 * 11 +  7] = 6'b001000;
assign fontdata[23 * 11 +  8] = 6'b001000;
assign fontdata[23 * 11 +  9] = 6'b000000;
assign fontdata[23 * 11 + 10] = 6'b000000;
assign fontdata[24 * 11 +  0] = 6'b000000;
assign fontdata[24 * 11 +  1] = 6'b000000;
assign fontdata[24 * 11 +  2] = 6'b011100;
assign fontdata[24 * 11 +  3] = 6'b100010;
assign fontdata[24 * 11 +  4] = 6'b100010;
assign fontdata[24 * 11 +  5] = 6'b011100;
assign fontdata[24 * 11 +  6] = 6'b100010;
assign fontdata[24 * 11 +  7] = 6'b100010;
assign fontdata[24 * 11 +  8] = 6'b011100;
assign fontdata[24 * 11 +  9] = 6'b000000;
assign fontdata[24 * 11 + 10] = 6'b000000;
assign fontdata[25 * 11 +  0] = 6'b000000;
assign fontdata[25 * 11 +  1] = 6'b000000;
assign fontdata[25 * 11 +  2] = 6'b011100;
assign fontdata[25 * 11 +  3] = 6'b100010;
assign fontdata[25 * 11 +  4] = 6'b100010;
assign fontdata[25 * 11 +  5] = 6'b011110;
assign fontdata[25 * 11 +  6] = 6'b000010;
assign fontdata[25 * 11 +  7] = 6'b000010;
assign fontdata[25 * 11 +  8] = 6'b011100;
assign fontdata[25 * 11 +  9] = 6'b000000;
assign fontdata[25 * 11 + 10] = 6'b000000;
assign fontdata[26 * 11 +  0] = 6'b000000;
assign fontdata[26 * 11 +  1] = 6'b000000;
assign fontdata[26 * 11 +  2] = 6'b000000;
assign fontdata[26 * 11 +  3] = 6'b000000;
assign fontdata[26 * 11 +  4] = 6'b001100;
assign fontdata[26 * 11 +  5] = 6'b001100;
assign fontdata[26 * 11 +  6] = 6'b000000;
assign fontdata[26 * 11 +  7] = 6'b001100;
assign fontdata[26 * 11 +  8] = 6'b001100;
assign fontdata[26 * 11 +  9] = 6'b000000;
assign fontdata[26 * 11 + 10] = 6'b000000;
assign fontdata[27 * 11 +  0] = 6'b000000;
assign fontdata[27 * 11 +  1] = 6'b000000;
assign fontdata[27 * 11 +  2] = 6'b000000;
assign fontdata[27 * 11 +  3] = 6'b000000;
assign fontdata[27 * 11 +  4] = 6'b011000;
assign fontdata[27 * 11 +  5] = 6'b011000;
assign fontdata[27 * 11 +  6] = 6'b000000;
assign fontdata[27 * 11 +  7] = 6'b011000;
assign fontdata[27 * 11 +  8] = 6'b011000;
assign fontdata[27 * 11 +  9] = 6'b001000;
assign fontdata[27 * 11 + 10] = 6'b010000;
assign fontdata[28 * 11 +  0] = 6'b000000;
assign fontdata[28 * 11 +  1] = 6'b000000;
assign fontdata[28 * 11 +  2] = 6'b000010;
assign fontdata[28 * 11 +  3] = 6'b000100;
assign fontdata[28 * 11 +  4] = 6'b001000;
assign fontdata[28 * 11 +  5] = 6'b010000;
assign fontdata[28 * 11 +  6] = 6'b001000;
assign fontdata[28 * 11 +  7] = 6'b000100;
assign fontdata[28 * 11 +  8] = 6'b000010;
assign fontdata[28 * 11 +  9] = 6'b000000;
assign fontdata[28 * 11 + 10] = 6'b000000;
assign fontdata[29 * 11 +  0] = 6'b000000;
assign fontdata[29 * 11 +  1] = 6'b000000;
assign fontdata[29 * 11 +  2] = 6'b000000;
assign fontdata[29 * 11 +  3] = 6'b000000;
assign fontdata[29 * 11 +  4] = 6'b111110;
assign fontdata[29 * 11 +  5] = 6'b000000;
assign fontdata[29 * 11 +  6] = 6'b111110;
assign fontdata[29 * 11 +  7] = 6'b000000;
assign fontdata[29 * 11 +  8] = 6'b000000;
assign fontdata[29 * 11 +  9] = 6'b000000;
assign fontdata[29 * 11 + 10] = 6'b000000;
assign fontdata[30 * 11 +  0] = 6'b000000;
assign fontdata[30 * 11 +  1] = 6'b000000;
assign fontdata[30 * 11 +  2] = 6'b010000;
assign fontdata[30 * 11 +  3] = 6'b001000;
assign fontdata[30 * 11 +  4] = 6'b000100;
assign fontdata[30 * 11 +  5] = 6'b000010;
assign fontdata[30 * 11 +  6] = 6'b000100;
assign fontdata[30 * 11 +  7] = 6'b001000;
assign fontdata[30 * 11 +  8] = 6'b010000;
assign fontdata[30 * 11 +  9] = 6'b000000;
assign fontdata[30 * 11 + 10] = 6'b000000;
assign fontdata[31 * 11 +  0] = 6'b000000;
assign fontdata[31 * 11 +  1] = 6'b000000;
assign fontdata[31 * 11 +  2] = 6'b011100;
assign fontdata[31 * 11 +  3] = 6'b100010;
assign fontdata[31 * 11 +  4] = 6'b000010;
assign fontdata[31 * 11 +  5] = 6'b000100;
assign fontdata[31 * 11 +  6] = 6'b001000;
assign fontdata[31 * 11 +  7] = 6'b000000;
assign fontdata[31 * 11 +  8] = 6'b001000;
assign fontdata[31 * 11 +  9] = 6'b000000;
assign fontdata[31 * 11 + 10] = 6'b000000;
assign fontdata[32 * 11 +  0] = 6'b000000;
assign fontdata[32 * 11 +  1] = 6'b000000;
assign fontdata[32 * 11 +  2] = 6'b011100;
assign fontdata[32 * 11 +  3] = 6'b100010;
assign fontdata[32 * 11 +  4] = 6'b101110;
assign fontdata[32 * 11 +  5] = 6'b101010;
assign fontdata[32 * 11 +  6] = 6'b101110;
assign fontdata[32 * 11 +  7] = 6'b100000;
assign fontdata[32 * 11 +  8] = 6'b011110;
assign fontdata[32 * 11 +  9] = 6'b000000;
assign fontdata[32 * 11 + 10] = 6'b000000;
assign fontdata[33 * 11 +  0] = 6'b000000;
assign fontdata[33 * 11 +  1] = 6'b011100;
assign fontdata[33 * 11 +  2] = 6'b100010;
assign fontdata[33 * 11 +  3] = 6'b100010;
assign fontdata[33 * 11 +  4] = 6'b111110;
assign fontdata[33 * 11 +  5] = 6'b100010;
assign fontdata[33 * 11 +  6] = 6'b100010;
assign fontdata[33 * 11 +  7] = 6'b100010;
assign fontdata[33 * 11 +  8] = 6'b100010;
assign fontdata[33 * 11 +  9] = 6'b000000;
assign fontdata[33 * 11 + 10] = 6'b000000;
assign fontdata[34 * 11 +  0] = 6'b000000;
assign fontdata[34 * 11 +  1] = 6'b111100;
assign fontdata[34 * 11 +  2] = 6'b100010;
assign fontdata[34 * 11 +  3] = 6'b100010;
assign fontdata[34 * 11 +  4] = 6'b111100;
assign fontdata[34 * 11 +  5] = 6'b100010;
assign fontdata[34 * 11 +  6] = 6'b100010;
assign fontdata[34 * 11 +  7] = 6'b100010;
assign fontdata[34 * 11 +  8] = 6'b111100;
assign fontdata[34 * 11 +  9] = 6'b000000;
assign fontdata[34 * 11 + 10] = 6'b000000;
assign fontdata[35 * 11 +  0] = 6'b000000;
assign fontdata[35 * 11 +  1] = 6'b011100;
assign fontdata[35 * 11 +  2] = 6'b100010;
assign fontdata[35 * 11 +  3] = 6'b100000;
assign fontdata[35 * 11 +  4] = 6'b100000;
assign fontdata[35 * 11 +  5] = 6'b100000;
assign fontdata[35 * 11 +  6] = 6'b100000;
assign fontdata[35 * 11 +  7] = 6'b100010;
assign fontdata[35 * 11 +  8] = 6'b011100;
assign fontdata[35 * 11 +  9] = 6'b000000;
assign fontdata[35 * 11 + 10] = 6'b000000;
assign fontdata[36 * 11 +  0] = 6'b000000;
assign fontdata[36 * 11 +  1] = 6'b111100;
assign fontdata[36 * 11 +  2] = 6'b100010;
assign fontdata[36 * 11 +  3] = 6'b100010;
assign fontdata[36 * 11 +  4] = 6'b100010;
assign fontdata[36 * 11 +  5] = 6'b100010;
assign fontdata[36 * 11 +  6] = 6'b100010;
assign fontdata[36 * 11 +  7] = 6'b100010;
assign fontdata[36 * 11 +  8] = 6'b111100;
assign fontdata[36 * 11 +  9] = 6'b000000;
assign fontdata[36 * 11 + 10] = 6'b000000;
assign fontdata[37 * 11 +  0] = 6'b000000;
assign fontdata[37 * 11 +  1] = 6'b111110;
assign fontdata[37 * 11 +  2] = 6'b100000;
assign fontdata[37 * 11 +  3] = 6'b100000;
assign fontdata[37 * 11 +  4] = 6'b111100;
assign fontdata[37 * 11 +  5] = 6'b100000;
assign fontdata[37 * 11 +  6] = 6'b100000;
assign fontdata[37 * 11 +  7] = 6'b100000;
assign fontdata[37 * 11 +  8] = 6'b111110;
assign fontdata[37 * 11 +  9] = 6'b000000;
assign fontdata[37 * 11 + 10] = 6'b000000;
assign fontdata[38 * 11 +  0] = 6'b000000;
assign fontdata[38 * 11 +  1] = 6'b111110;
assign fontdata[38 * 11 +  2] = 6'b100000;
assign fontdata[38 * 11 +  3] = 6'b100000;
assign fontdata[38 * 11 +  4] = 6'b111100;
assign fontdata[38 * 11 +  5] = 6'b100000;
assign fontdata[38 * 11 +  6] = 6'b100000;
assign fontdata[38 * 11 +  7] = 6'b100000;
assign fontdata[38 * 11 +  8] = 6'b100000;
assign fontdata[38 * 11 +  9] = 6'b000000;
assign fontdata[38 * 11 + 10] = 6'b000000;
assign fontdata[39 * 11 +  0] = 6'b000000;
assign fontdata[39 * 11 +  1] = 6'b011100;
assign fontdata[39 * 11 +  2] = 6'b100010;
assign fontdata[39 * 11 +  3] = 6'b100000;
assign fontdata[39 * 11 +  4] = 6'b101110;
assign fontdata[39 * 11 +  5] = 6'b100010;
assign fontdata[39 * 11 +  6] = 6'b100010;
assign fontdata[39 * 11 +  7] = 6'b100010;
assign fontdata[39 * 11 +  8] = 6'b011100;
assign fontdata[39 * 11 +  9] = 6'b000000;
assign fontdata[39 * 11 + 10] = 6'b000000;
assign fontdata[40 * 11 +  0] = 6'b000000;
assign fontdata[40 * 11 +  1] = 6'b100010;
assign fontdata[40 * 11 +  2] = 6'b100010;
assign fontdata[40 * 11 +  3] = 6'b100010;
assign fontdata[40 * 11 +  4] = 6'b111110;
assign fontdata[40 * 11 +  5] = 6'b100010;
assign fontdata[40 * 11 +  6] = 6'b100010;
assign fontdata[40 * 11 +  7] = 6'b100010;
assign fontdata[40 * 11 +  8] = 6'b100010;
assign fontdata[40 * 11 +  9] = 6'b000000;
assign fontdata[40 * 11 + 10] = 6'b000000;
assign fontdata[41 * 11 +  0] = 6'b000000;
assign fontdata[41 * 11 +  1] = 6'b011100;
assign fontdata[41 * 11 +  2] = 6'b001000;
assign fontdata[41 * 11 +  3] = 6'b001000;
assign fontdata[41 * 11 +  4] = 6'b001000;
assign fontdata[41 * 11 +  5] = 6'b001000;
assign fontdata[41 * 11 +  6] = 6'b001000;
assign fontdata[41 * 11 +  7] = 6'b001000;
assign fontdata[41 * 11 +  8] = 6'b011100;
assign fontdata[41 * 11 +  9] = 6'b000000;
assign fontdata[41 * 11 + 10] = 6'b000000;
assign fontdata[42 * 11 +  0] = 6'b000000;
assign fontdata[42 * 11 +  1] = 6'b000010;
assign fontdata[42 * 11 +  2] = 6'b000010;
assign fontdata[42 * 11 +  3] = 6'b000010;
assign fontdata[42 * 11 +  4] = 6'b000010;
assign fontdata[42 * 11 +  5] = 6'b000010;
assign fontdata[42 * 11 +  6] = 6'b100010;
assign fontdata[42 * 11 +  7] = 6'b100010;
assign fontdata[42 * 11 +  8] = 6'b011100;
assign fontdata[42 * 11 +  9] = 6'b000000;
assign fontdata[42 * 11 + 10] = 6'b000000;
assign fontdata[43 * 11 +  0] = 6'b000000;
assign fontdata[43 * 11 +  1] = 6'b100010;
assign fontdata[43 * 11 +  2] = 6'b100100;
assign fontdata[43 * 11 +  3] = 6'b101000;
assign fontdata[43 * 11 +  4] = 6'b110000;
assign fontdata[43 * 11 +  5] = 6'b101000;
assign fontdata[43 * 11 +  6] = 6'b100100;
assign fontdata[43 * 11 +  7] = 6'b100010;
assign fontdata[43 * 11 +  8] = 6'b100010;
assign fontdata[43 * 11 +  9] = 6'b000000;
assign fontdata[43 * 11 + 10] = 6'b000000;
assign fontdata[44 * 11 +  0] = 6'b000000;
assign fontdata[44 * 11 +  1] = 6'b100000;
assign fontdata[44 * 11 +  2] = 6'b100000;
assign fontdata[44 * 11 +  3] = 6'b100000;
assign fontdata[44 * 11 +  4] = 6'b100000;
assign fontdata[44 * 11 +  5] = 6'b100000;
assign fontdata[44 * 11 +  6] = 6'b100000;
assign fontdata[44 * 11 +  7] = 6'b100000;
assign fontdata[44 * 11 +  8] = 6'b111110;
assign fontdata[44 * 11 +  9] = 6'b000000;
assign fontdata[44 * 11 + 10] = 6'b000000;
assign fontdata[45 * 11 +  0] = 6'b000000;
assign fontdata[45 * 11 +  1] = 6'b100010;
assign fontdata[45 * 11 +  2] = 6'b110110;
assign fontdata[45 * 11 +  3] = 6'b101010;
assign fontdata[45 * 11 +  4] = 6'b101010;
assign fontdata[45 * 11 +  5] = 6'b100010;
assign fontdata[45 * 11 +  6] = 6'b100010;
assign fontdata[45 * 11 +  7] = 6'b100010;
assign fontdata[45 * 11 +  8] = 6'b100010;
assign fontdata[45 * 11 +  9] = 6'b000000;
assign fontdata[45 * 11 + 10] = 6'b000000;
assign fontdata[46 * 11 +  0] = 6'b000000;
assign fontdata[46 * 11 +  1] = 6'b100010;
assign fontdata[46 * 11 +  2] = 6'b110010;
assign fontdata[46 * 11 +  3] = 6'b110010;
assign fontdata[46 * 11 +  4] = 6'b101010;
assign fontdata[46 * 11 +  5] = 6'b101010;
assign fontdata[46 * 11 +  6] = 6'b100110;
assign fontdata[46 * 11 +  7] = 6'b100110;
assign fontdata[46 * 11 +  8] = 6'b100010;
assign fontdata[46 * 11 +  9] = 6'b000000;
assign fontdata[46 * 11 + 10] = 6'b000000;
assign fontdata[47 * 11 +  0] = 6'b000000;
assign fontdata[47 * 11 +  1] = 6'b011100;
assign fontdata[47 * 11 +  2] = 6'b100010;
assign fontdata[47 * 11 +  3] = 6'b100010;
assign fontdata[47 * 11 +  4] = 6'b100010;
assign fontdata[47 * 11 +  5] = 6'b100010;
assign fontdata[47 * 11 +  6] = 6'b100010;
assign fontdata[47 * 11 +  7] = 6'b100010;
assign fontdata[47 * 11 +  8] = 6'b011100;
assign fontdata[47 * 11 +  9] = 6'b000000;
assign fontdata[47 * 11 + 10] = 6'b000000;
assign fontdata[48 * 11 +  0] = 6'b000000;
assign fontdata[48 * 11 +  1] = 6'b111100;
assign fontdata[48 * 11 +  2] = 6'b100010;
assign fontdata[48 * 11 +  3] = 6'b100010;
assign fontdata[48 * 11 +  4] = 6'b111100;
assign fontdata[48 * 11 +  5] = 6'b100000;
assign fontdata[48 * 11 +  6] = 6'b100000;
assign fontdata[48 * 11 +  7] = 6'b100000;
assign fontdata[48 * 11 +  8] = 6'b100000;
assign fontdata[48 * 11 +  9] = 6'b000000;
assign fontdata[48 * 11 + 10] = 6'b000000;
assign fontdata[49 * 11 +  0] = 6'b000000;
assign fontdata[49 * 11 +  1] = 6'b011100;
assign fontdata[49 * 11 +  2] = 6'b100010;
assign fontdata[49 * 11 +  3] = 6'b100010;
assign fontdata[49 * 11 +  4] = 6'b100010;
assign fontdata[49 * 11 +  5] = 6'b100010;
assign fontdata[49 * 11 +  6] = 6'b101010;
assign fontdata[49 * 11 +  7] = 6'b100100;
assign fontdata[49 * 11 +  8] = 6'b011010;
assign fontdata[49 * 11 +  9] = 6'b000010;
assign fontdata[49 * 11 + 10] = 6'b000000;
assign fontdata[50 * 11 +  0] = 6'b000000;
assign fontdata[50 * 11 +  1] = 6'b111100;
assign fontdata[50 * 11 +  2] = 6'b100010;
assign fontdata[50 * 11 +  3] = 6'b100010;
assign fontdata[50 * 11 +  4] = 6'b111100;
assign fontdata[50 * 11 +  5] = 6'b100100;
assign fontdata[50 * 11 +  6] = 6'b100010;
assign fontdata[50 * 11 +  7] = 6'b100010;
assign fontdata[50 * 11 +  8] = 6'b100010;
assign fontdata[50 * 11 +  9] = 6'b000000;
assign fontdata[50 * 11 + 10] = 6'b000000;
assign fontdata[51 * 11 +  0] = 6'b000000;
assign fontdata[51 * 11 +  1] = 6'b011100;
assign fontdata[51 * 11 +  2] = 6'b100010;
assign fontdata[51 * 11 +  3] = 6'b100000;
assign fontdata[51 * 11 +  4] = 6'b011100;
assign fontdata[51 * 11 +  5] = 6'b000010;
assign fontdata[51 * 11 +  6] = 6'b000010;
assign fontdata[51 * 11 +  7] = 6'b100010;
assign fontdata[51 * 11 +  8] = 6'b011100;
assign fontdata[51 * 11 +  9] = 6'b000000;
assign fontdata[51 * 11 + 10] = 6'b000000;
assign fontdata[52 * 11 +  0] = 6'b000000;
assign fontdata[52 * 11 +  1] = 6'b111110;
assign fontdata[52 * 11 +  2] = 6'b001000;
assign fontdata[52 * 11 +  3] = 6'b001000;
assign fontdata[52 * 11 +  4] = 6'b001000;
assign fontdata[52 * 11 +  5] = 6'b001000;
assign fontdata[52 * 11 +  6] = 6'b001000;
assign fontdata[52 * 11 +  7] = 6'b001000;
assign fontdata[52 * 11 +  8] = 6'b001000;
assign fontdata[52 * 11 +  9] = 6'b000000;
assign fontdata[52 * 11 + 10] = 6'b000000;
assign fontdata[53 * 11 +  0] = 6'b000000;
assign fontdata[53 * 11 +  1] = 6'b100010;
assign fontdata[53 * 11 +  2] = 6'b100010;
assign fontdata[53 * 11 +  3] = 6'b100010;
assign fontdata[53 * 11 +  4] = 6'b100010;
assign fontdata[53 * 11 +  5] = 6'b100010;
assign fontdata[53 * 11 +  6] = 6'b100010;
assign fontdata[53 * 11 +  7] = 6'b100010;
assign fontdata[53 * 11 +  8] = 6'b011100;
assign fontdata[53 * 11 +  9] = 6'b000000;
assign fontdata[53 * 11 + 10] = 6'b000000;
assign fontdata[54 * 11 +  0] = 6'b000000;
assign fontdata[54 * 11 +  1] = 6'b100010;
assign fontdata[54 * 11 +  2] = 6'b100010;
assign fontdata[54 * 11 +  3] = 6'b100010;
assign fontdata[54 * 11 +  4] = 6'b100010;
assign fontdata[54 * 11 +  5] = 6'b010100;
assign fontdata[54 * 11 +  6] = 6'b010100;
assign fontdata[54 * 11 +  7] = 6'b001000;
assign fontdata[54 * 11 +  8] = 6'b001000;
assign fontdata[54 * 11 +  9] = 6'b000000;
assign fontdata[54 * 11 + 10] = 6'b000000;
assign fontdata[55 * 11 +  0] = 6'b000000;
assign fontdata[55 * 11 +  1] = 6'b100010;
assign fontdata[55 * 11 +  2] = 6'b100010;
assign fontdata[55 * 11 +  3] = 6'b100010;
assign fontdata[55 * 11 +  4] = 6'b101010;
assign fontdata[55 * 11 +  5] = 6'b101010;
assign fontdata[55 * 11 +  6] = 6'b101010;
assign fontdata[55 * 11 +  7] = 6'b010100;
assign fontdata[55 * 11 +  8] = 6'b010100;
assign fontdata[55 * 11 +  9] = 6'b000000;
assign fontdata[55 * 11 + 10] = 6'b000000;
assign fontdata[56 * 11 +  0] = 6'b000000;
assign fontdata[56 * 11 +  1] = 6'b100010;
assign fontdata[56 * 11 +  2] = 6'b100010;
assign fontdata[56 * 11 +  3] = 6'b010100;
assign fontdata[56 * 11 +  4] = 6'b001000;
assign fontdata[56 * 11 +  5] = 6'b010100;
assign fontdata[56 * 11 +  6] = 6'b100010;
assign fontdata[56 * 11 +  7] = 6'b100010;
assign fontdata[56 * 11 +  8] = 6'b100010;
assign fontdata[56 * 11 +  9] = 6'b000000;
assign fontdata[56 * 11 + 10] = 6'b000000;
assign fontdata[57 * 11 +  0] = 6'b000000;
assign fontdata[57 * 11 +  1] = 6'b100010;
assign fontdata[57 * 11 +  2] = 6'b100010;
assign fontdata[57 * 11 +  3] = 6'b010100;
assign fontdata[57 * 11 +  4] = 6'b001000;
assign fontdata[57 * 11 +  5] = 6'b001000;
assign fontdata[57 * 11 +  6] = 6'b001000;
assign fontdata[57 * 11 +  7] = 6'b001000;
assign fontdata[57 * 11 +  8] = 6'b001000;
assign fontdata[57 * 11 +  9] = 6'b000000;
assign fontdata[57 * 11 + 10] = 6'b000000;
assign fontdata[58 * 11 +  0] = 6'b000000;
assign fontdata[58 * 11 +  1] = 6'b111110;
assign fontdata[58 * 11 +  2] = 6'b000010;
assign fontdata[58 * 11 +  3] = 6'b000100;
assign fontdata[58 * 11 +  4] = 6'b001000;
assign fontdata[58 * 11 +  5] = 6'b010000;
assign fontdata[58 * 11 +  6] = 6'b100000;
assign fontdata[58 * 11 +  7] = 6'b100000;
assign fontdata[58 * 11 +  8] = 6'b111110;
assign fontdata[58 * 11 +  9] = 6'b000000;
assign fontdata[58 * 11 + 10] = 6'b000000;
assign fontdata[59 * 11 +  0] = 6'b000000;
assign fontdata[59 * 11 +  1] = 6'b001110;
assign fontdata[59 * 11 +  2] = 6'b001000;
assign fontdata[59 * 11 +  3] = 6'b001000;
assign fontdata[59 * 11 +  4] = 6'b001000;
assign fontdata[59 * 11 +  5] = 6'b001000;
assign fontdata[59 * 11 +  6] = 6'b001000;
assign fontdata[59 * 11 +  7] = 6'b001000;
assign fontdata[59 * 11 +  8] = 6'b001000;
assign fontdata[59 * 11 +  9] = 6'b001110;
assign fontdata[59 * 11 + 10] = 6'b000000;
assign fontdata[60 * 11 +  0] = 6'b000000;
assign fontdata[60 * 11 +  1] = 6'b010000;
assign fontdata[60 * 11 +  2] = 6'b010000;
assign fontdata[60 * 11 +  3] = 6'b001000;
assign fontdata[60 * 11 +  4] = 6'b001000;
assign fontdata[60 * 11 +  5] = 6'b000100;
assign fontdata[60 * 11 +  6] = 6'b000100;
assign fontdata[60 * 11 +  7] = 6'b000010;
assign fontdata[60 * 11 +  8] = 6'b000010;
assign fontdata[60 * 11 +  9] = 6'b000001;
assign fontdata[60 * 11 + 10] = 6'b000001;
assign fontdata[61 * 11 +  0] = 6'b000000;
assign fontdata[61 * 11 +  1] = 6'b111000;
assign fontdata[61 * 11 +  2] = 6'b001000;
assign fontdata[61 * 11 +  3] = 6'b001000;
assign fontdata[61 * 11 +  4] = 6'b001000;
assign fontdata[61 * 11 +  5] = 6'b001000;
assign fontdata[61 * 11 +  6] = 6'b001000;
assign fontdata[61 * 11 +  7] = 6'b001000;
assign fontdata[61 * 11 +  8] = 6'b001000;
assign fontdata[61 * 11 +  9] = 6'b111000;
assign fontdata[61 * 11 + 10] = 6'b000000;
assign fontdata[62 * 11 +  0] = 6'b000000;
assign fontdata[62 * 11 +  1] = 6'b000000;
assign fontdata[62 * 11 +  2] = 6'b001000;
assign fontdata[62 * 11 +  3] = 6'b010100;
assign fontdata[62 * 11 +  4] = 6'b100010;
assign fontdata[62 * 11 +  5] = 6'b000000;
assign fontdata[62 * 11 +  6] = 6'b000000;
assign fontdata[62 * 11 +  7] = 6'b000000;
assign fontdata[62 * 11 +  8] = 6'b000000;
assign fontdata[62 * 11 +  9] = 6'b000000;
assign fontdata[62 * 11 + 10] = 6'b000000;
assign fontdata[63 * 11 +  0] = 6'b000000;
assign fontdata[63 * 11 +  1] = 6'b000000;
assign fontdata[63 * 11 +  2] = 6'b000000;
assign fontdata[63 * 11 +  3] = 6'b000000;
assign fontdata[63 * 11 +  4] = 6'b000000;
assign fontdata[63 * 11 +  5] = 6'b000000;
assign fontdata[63 * 11 +  6] = 6'b000000;
assign fontdata[63 * 11 +  7] = 6'b000000;
assign fontdata[63 * 11 +  8] = 6'b000000;
assign fontdata[63 * 11 +  9] = 6'b111111;
assign fontdata[63 * 11 + 10] = 6'b000000;
assign fontdata[64 * 11 +  0] = 6'b000000;
assign fontdata[64 * 11 +  1] = 6'b010000;
assign fontdata[64 * 11 +  2] = 6'b001000;
assign fontdata[64 * 11 +  3] = 6'b000100;
assign fontdata[64 * 11 +  4] = 6'b000000;
assign fontdata[64 * 11 +  5] = 6'b000000;
assign fontdata[64 * 11 +  6] = 6'b000000;
assign fontdata[64 * 11 +  7] = 6'b000000;
assign fontdata[64 * 11 +  8] = 6'b000000;
assign fontdata[64 * 11 +  9] = 6'b000000;
assign fontdata[64 * 11 + 10] = 6'b000000;
assign fontdata[65 * 11 +  0] = 6'b000000;
assign fontdata[65 * 11 +  1] = 6'b000000;
assign fontdata[65 * 11 +  2] = 6'b000000;
assign fontdata[65 * 11 +  3] = 6'b000000;
assign fontdata[65 * 11 +  4] = 6'b011100;
assign fontdata[65 * 11 +  5] = 6'b000010;
assign fontdata[65 * 11 +  6] = 6'b011110;
assign fontdata[65 * 11 +  7] = 6'b100010;
assign fontdata[65 * 11 +  8] = 6'b011110;
assign fontdata[65 * 11 +  9] = 6'b000000;
assign fontdata[65 * 11 + 10] = 6'b000000;
assign fontdata[66 * 11 +  0] = 6'b000000;
assign fontdata[66 * 11 +  1] = 6'b100000;
assign fontdata[66 * 11 +  2] = 6'b100000;
assign fontdata[66 * 11 +  3] = 6'b100000;
assign fontdata[66 * 11 +  4] = 6'b101100;
assign fontdata[66 * 11 +  5] = 6'b110010;
assign fontdata[66 * 11 +  6] = 6'b100010;
assign fontdata[66 * 11 +  7] = 6'b100010;
assign fontdata[66 * 11 +  8] = 6'b111100;
assign fontdata[66 * 11 +  9] = 6'b000000;
assign fontdata[66 * 11 + 10] = 6'b000000;
assign fontdata[67 * 11 +  0] = 6'b000000;
assign fontdata[67 * 11 +  1] = 6'b000000;
assign fontdata[67 * 11 +  2] = 6'b000000;
assign fontdata[67 * 11 +  3] = 6'b000000;
assign fontdata[67 * 11 +  4] = 6'b011110;
assign fontdata[67 * 11 +  5] = 6'b100000;
assign fontdata[67 * 11 +  6] = 6'b100000;
assign fontdata[67 * 11 +  7] = 6'b100000;
assign fontdata[67 * 11 +  8] = 6'b011110;
assign fontdata[67 * 11 +  9] = 6'b000000;
assign fontdata[67 * 11 + 10] = 6'b000000;
assign fontdata[68 * 11 +  0] = 6'b000000;
assign fontdata[68 * 11 +  1] = 6'b000010;
assign fontdata[68 * 11 +  2] = 6'b000010;
assign fontdata[68 * 11 +  3] = 6'b000010;
assign fontdata[68 * 11 +  4] = 6'b011110;
assign fontdata[68 * 11 +  5] = 6'b100010;
assign fontdata[68 * 11 +  6] = 6'b100010;
assign fontdata[68 * 11 +  7] = 6'b100110;
assign fontdata[68 * 11 +  8] = 6'b011010;
assign fontdata[68 * 11 +  9] = 6'b000000;
assign fontdata[68 * 11 + 10] = 6'b000000;
assign fontdata[69 * 11 +  0] = 6'b000000;
assign fontdata[69 * 11 +  1] = 6'b000000;
assign fontdata[69 * 11 +  2] = 6'b000000;
assign fontdata[69 * 11 +  3] = 6'b000000;
assign fontdata[69 * 11 +  4] = 6'b011100;
assign fontdata[69 * 11 +  5] = 6'b100010;
assign fontdata[69 * 11 +  6] = 6'b111110;
assign fontdata[69 * 11 +  7] = 6'b100000;
assign fontdata[69 * 11 +  8] = 6'b011110;
assign fontdata[69 * 11 +  9] = 6'b000000;
assign fontdata[69 * 11 + 10] = 6'b000000;
assign fontdata[70 * 11 +  0] = 6'b000000;
assign fontdata[70 * 11 +  1] = 6'b001100;
assign fontdata[70 * 11 +  2] = 6'b010000;
assign fontdata[70 * 11 +  3] = 6'b010000;
assign fontdata[70 * 11 +  4] = 6'b011100;
assign fontdata[70 * 11 +  5] = 6'b010000;
assign fontdata[70 * 11 +  6] = 6'b010000;
assign fontdata[70 * 11 +  7] = 6'b010000;
assign fontdata[70 * 11 +  8] = 6'b010000;
assign fontdata[70 * 11 +  9] = 6'b000000;
assign fontdata[70 * 11 + 10] = 6'b000000;
assign fontdata[71 * 11 +  0] = 6'b000000;
assign fontdata[71 * 11 +  1] = 6'b000000;
assign fontdata[71 * 11 +  2] = 6'b000000;
assign fontdata[71 * 11 +  3] = 6'b000000;
assign fontdata[71 * 11 +  4] = 6'b011110;
assign fontdata[71 * 11 +  5] = 6'b100010;
assign fontdata[71 * 11 +  6] = 6'b100010;
assign fontdata[71 * 11 +  7] = 6'b100110;
assign fontdata[71 * 11 +  8] = 6'b011010;
assign fontdata[71 * 11 +  9] = 6'b000010;
assign fontdata[71 * 11 + 10] = 6'b011100;
assign fontdata[72 * 11 +  0] = 6'b000000;
assign fontdata[72 * 11 +  1] = 6'b100000;
assign fontdata[72 * 11 +  2] = 6'b100000;
assign fontdata[72 * 11 +  3] = 6'b100000;
assign fontdata[72 * 11 +  4] = 6'b101100;
assign fontdata[72 * 11 +  5] = 6'b110010;
assign fontdata[72 * 11 +  6] = 6'b100010;
assign fontdata[72 * 11 +  7] = 6'b100010;
assign fontdata[72 * 11 +  8] = 6'b100010;
assign fontdata[72 * 11 +  9] = 6'b000000;
assign fontdata[72 * 11 + 10] = 6'b000000;
assign fontdata[73 * 11 +  0] = 6'b000000;
assign fontdata[73 * 11 +  1] = 6'b000000;
assign fontdata[73 * 11 +  2] = 6'b001000;
assign fontdata[73 * 11 +  3] = 6'b000000;
assign fontdata[73 * 11 +  4] = 6'b011000;
assign fontdata[73 * 11 +  5] = 6'b001000;
assign fontdata[73 * 11 +  6] = 6'b001000;
assign fontdata[73 * 11 +  7] = 6'b001000;
assign fontdata[73 * 11 +  8] = 6'b001100;
assign fontdata[73 * 11 +  9] = 6'b000000;
assign fontdata[73 * 11 + 10] = 6'b000000;
assign fontdata[74 * 11 +  0] = 6'b000000;
assign fontdata[74 * 11 +  1] = 6'b000000;
assign fontdata[74 * 11 +  2] = 6'b001000;
assign fontdata[74 * 11 +  3] = 6'b000000;
assign fontdata[74 * 11 +  4] = 6'b011000;
assign fontdata[74 * 11 +  5] = 6'b001000;
assign fontdata[74 * 11 +  6] = 6'b001000;
assign fontdata[74 * 11 +  7] = 6'b001000;
assign fontdata[74 * 11 +  8] = 6'b001000;
assign fontdata[74 * 11 +  9] = 6'b001000;
assign fontdata[74 * 11 + 10] = 6'b110000;
assign fontdata[75 * 11 +  0] = 6'b000000;
assign fontdata[75 * 11 +  1] = 6'b100000;
assign fontdata[75 * 11 +  2] = 6'b100000;
assign fontdata[75 * 11 +  3] = 6'b100000;
assign fontdata[75 * 11 +  4] = 6'b100100;
assign fontdata[75 * 11 +  5] = 6'b101000;
assign fontdata[75 * 11 +  6] = 6'b111000;
assign fontdata[75 * 11 +  7] = 6'b100100;
assign fontdata[75 * 11 +  8] = 6'b100010;
assign fontdata[75 * 11 +  9] = 6'b000000;
assign fontdata[75 * 11 + 10] = 6'b000000;
assign fontdata[76 * 11 +  0] = 6'b000000;
assign fontdata[76 * 11 +  1] = 6'b011000;
assign fontdata[76 * 11 +  2] = 6'b001000;
assign fontdata[76 * 11 +  3] = 6'b001000;
assign fontdata[76 * 11 +  4] = 6'b001000;
assign fontdata[76 * 11 +  5] = 6'b001000;
assign fontdata[76 * 11 +  6] = 6'b001000;
assign fontdata[76 * 11 +  7] = 6'b001000;
assign fontdata[76 * 11 +  8] = 6'b000110;
assign fontdata[76 * 11 +  9] = 6'b000000;
assign fontdata[76 * 11 + 10] = 6'b000000;
assign fontdata[77 * 11 +  0] = 6'b000000;
assign fontdata[77 * 11 +  1] = 6'b000000;
assign fontdata[77 * 11 +  2] = 6'b000000;
assign fontdata[77 * 11 +  3] = 6'b000000;
assign fontdata[77 * 11 +  4] = 6'b111100;
assign fontdata[77 * 11 +  5] = 6'b101010;
assign fontdata[77 * 11 +  6] = 6'b101010;
assign fontdata[77 * 11 +  7] = 6'b101010;
assign fontdata[77 * 11 +  8] = 6'b101010;
assign fontdata[77 * 11 +  9] = 6'b000000;
assign fontdata[77 * 11 + 10] = 6'b000000;
assign fontdata[78 * 11 +  0] = 6'b000000;
assign fontdata[78 * 11 +  1] = 6'b000000;
assign fontdata[78 * 11 +  2] = 6'b000000;
assign fontdata[78 * 11 +  3] = 6'b000000;
assign fontdata[78 * 11 +  4] = 6'b111100;
assign fontdata[78 * 11 +  5] = 6'b100010;
assign fontdata[78 * 11 +  6] = 6'b100010;
assign fontdata[78 * 11 +  7] = 6'b100010;
assign fontdata[78 * 11 +  8] = 6'b100010;
assign fontdata[78 * 11 +  9] = 6'b000000;
assign fontdata[78 * 11 + 10] = 6'b000000;
assign fontdata[79 * 11 +  0] = 6'b000000;
assign fontdata[79 * 11 +  1] = 6'b000000;
assign fontdata[79 * 11 +  2] = 6'b000000;
assign fontdata[79 * 11 +  3] = 6'b000000;
assign fontdata[79 * 11 +  4] = 6'b011100;
assign fontdata[79 * 11 +  5] = 6'b100010;
assign fontdata[79 * 11 +  6] = 6'b100010;
assign fontdata[79 * 11 +  7] = 6'b100010;
assign fontdata[79 * 11 +  8] = 6'b011100;
assign fontdata[79 * 11 +  9] = 6'b000000;
assign fontdata[79 * 11 + 10] = 6'b000000;
assign fontdata[80 * 11 +  0] = 6'b000000;
assign fontdata[80 * 11 +  1] = 6'b000000;
assign fontdata[80 * 11 +  2] = 6'b000000;
assign fontdata[80 * 11 +  3] = 6'b000000;
assign fontdata[80 * 11 +  4] = 6'b101100;
assign fontdata[80 * 11 +  5] = 6'b110010;
assign fontdata[80 * 11 +  6] = 6'b100010;
assign fontdata[80 * 11 +  7] = 6'b100010;
assign fontdata[80 * 11 +  8] = 6'b111100;
assign fontdata[80 * 11 +  9] = 6'b100000;
assign fontdata[80 * 11 + 10] = 6'b100000;
assign fontdata[81 * 11 +  0] = 6'b000000;
assign fontdata[81 * 11 +  1] = 6'b000000;
assign fontdata[81 * 11 +  2] = 6'b000000;
assign fontdata[81 * 11 +  3] = 6'b000000;
assign fontdata[81 * 11 +  4] = 6'b011110;
assign fontdata[81 * 11 +  5] = 6'b100010;
assign fontdata[81 * 11 +  6] = 6'b100010;
assign fontdata[81 * 11 +  7] = 6'b100110;
assign fontdata[81 * 11 +  8] = 6'b011010;
assign fontdata[81 * 11 +  9] = 6'b000010;
assign fontdata[81 * 11 + 10] = 6'b000010;
assign fontdata[82 * 11 +  0] = 6'b000000;
assign fontdata[82 * 11 +  1] = 6'b000000;
assign fontdata[82 * 11 +  2] = 6'b000000;
assign fontdata[82 * 11 +  3] = 6'b000000;
assign fontdata[82 * 11 +  4] = 6'b101100;
assign fontdata[82 * 11 +  5] = 6'b110010;
assign fontdata[82 * 11 +  6] = 6'b100000;
assign fontdata[82 * 11 +  7] = 6'b100000;
assign fontdata[82 * 11 +  8] = 6'b100000;
assign fontdata[82 * 11 +  9] = 6'b000000;
assign fontdata[82 * 11 + 10] = 6'b000000;
assign fontdata[83 * 11 +  0] = 6'b000000;
assign fontdata[83 * 11 +  1] = 6'b000000;
assign fontdata[83 * 11 +  2] = 6'b000000;
assign fontdata[83 * 11 +  3] = 6'b000000;
assign fontdata[83 * 11 +  4] = 6'b011100;
assign fontdata[83 * 11 +  5] = 6'b100000;
assign fontdata[83 * 11 +  6] = 6'b011100;
assign fontdata[83 * 11 +  7] = 6'b000010;
assign fontdata[83 * 11 +  8] = 6'b111100;
assign fontdata[83 * 11 +  9] = 6'b000000;
assign fontdata[83 * 11 + 10] = 6'b000000;
assign fontdata[84 * 11 +  0] = 6'b000000;
assign fontdata[84 * 11 +  1] = 6'b010000;
assign fontdata[84 * 11 +  2] = 6'b010000;
assign fontdata[84 * 11 +  3] = 6'b010000;
assign fontdata[84 * 11 +  4] = 6'b111100;
assign fontdata[84 * 11 +  5] = 6'b010000;
assign fontdata[84 * 11 +  6] = 6'b010000;
assign fontdata[84 * 11 +  7] = 6'b010000;
assign fontdata[84 * 11 +  8] = 6'b001100;
assign fontdata[84 * 11 +  9] = 6'b000000;
assign fontdata[84 * 11 + 10] = 6'b000000;
assign fontdata[85 * 11 +  0] = 6'b000000;
assign fontdata[85 * 11 +  1] = 6'b000000;
assign fontdata[85 * 11 +  2] = 6'b000000;
assign fontdata[85 * 11 +  3] = 6'b000000;
assign fontdata[85 * 11 +  4] = 6'b100010;
assign fontdata[85 * 11 +  5] = 6'b100010;
assign fontdata[85 * 11 +  6] = 6'b100010;
assign fontdata[85 * 11 +  7] = 6'b100110;
assign fontdata[85 * 11 +  8] = 6'b011010;
assign fontdata[85 * 11 +  9] = 6'b000000;
assign fontdata[85 * 11 + 10] = 6'b000000;
assign fontdata[86 * 11 +  0] = 6'b000000;
assign fontdata[86 * 11 +  1] = 6'b000000;
assign fontdata[86 * 11 +  2] = 6'b000000;
assign fontdata[86 * 11 +  3] = 6'b000000;
assign fontdata[86 * 11 +  4] = 6'b100010;
assign fontdata[86 * 11 +  5] = 6'b100010;
assign fontdata[86 * 11 +  6] = 6'b010100;
assign fontdata[86 * 11 +  7] = 6'b010100;
assign fontdata[86 * 11 +  8] = 6'b001000;
assign fontdata[86 * 11 +  9] = 6'b000000;
assign fontdata[86 * 11 + 10] = 6'b000000;
assign fontdata[87 * 11 +  0] = 6'b000000;
assign fontdata[87 * 11 +  1] = 6'b000000;
assign fontdata[87 * 11 +  2] = 6'b000000;
assign fontdata[87 * 11 +  3] = 6'b000000;
assign fontdata[87 * 11 +  4] = 6'b100010;
assign fontdata[87 * 11 +  5] = 6'b101010;
assign fontdata[87 * 11 +  6] = 6'b101010;
assign fontdata[87 * 11 +  7] = 6'b101010;
assign fontdata[87 * 11 +  8] = 6'b010100;
assign fontdata[87 * 11 +  9] = 6'b000000;
assign fontdata[87 * 11 + 10] = 6'b000000;
assign fontdata[88 * 11 +  0] = 6'b000000;
assign fontdata[88 * 11 +  1] = 6'b000000;
assign fontdata[88 * 11 +  2] = 6'b000000;
assign fontdata[88 * 11 +  3] = 6'b000000;
assign fontdata[88 * 11 +  4] = 6'b100010;
assign fontdata[88 * 11 +  5] = 6'b010100;
assign fontdata[88 * 11 +  6] = 6'b001000;
assign fontdata[88 * 11 +  7] = 6'b010100;
assign fontdata[88 * 11 +  8] = 6'b100010;
assign fontdata[88 * 11 +  9] = 6'b000000;
assign fontdata[88 * 11 + 10] = 6'b000000;
assign fontdata[89 * 11 +  0] = 6'b000000;
assign fontdata[89 * 11 +  1] = 6'b000000;
assign fontdata[89 * 11 +  2] = 6'b000000;
assign fontdata[89 * 11 +  3] = 6'b000000;
assign fontdata[89 * 11 +  4] = 6'b100010;
assign fontdata[89 * 11 +  5] = 6'b100010;
assign fontdata[89 * 11 +  6] = 6'b100010;
assign fontdata[89 * 11 +  7] = 6'b100110;
assign fontdata[89 * 11 +  8] = 6'b011010;
assign fontdata[89 * 11 +  9] = 6'b000010;
assign fontdata[89 * 11 + 10] = 6'b011100;
assign fontdata[90 * 11 +  0] = 6'b000000;
assign fontdata[90 * 11 +  1] = 6'b000000;
assign fontdata[90 * 11 +  2] = 6'b000000;
assign fontdata[90 * 11 +  3] = 6'b000000;
assign fontdata[90 * 11 +  4] = 6'b111110;
assign fontdata[90 * 11 +  5] = 6'b000100;
assign fontdata[90 * 11 +  6] = 6'b001000;
assign fontdata[90 * 11 +  7] = 6'b010000;
assign fontdata[90 * 11 +  8] = 6'b111110;
assign fontdata[90 * 11 +  9] = 6'b000000;
assign fontdata[90 * 11 + 10] = 6'b000000;
assign fontdata[91 * 11 +  0] = 6'b000110;
assign fontdata[91 * 11 +  1] = 6'b001000;
assign fontdata[91 * 11 +  2] = 6'b001000;
assign fontdata[91 * 11 +  3] = 6'b001000;
assign fontdata[91 * 11 +  4] = 6'b001000;
assign fontdata[91 * 11 +  5] = 6'b110000;
assign fontdata[91 * 11 +  6] = 6'b001000;
assign fontdata[91 * 11 +  7] = 6'b001000;
assign fontdata[91 * 11 +  8] = 6'b001000;
assign fontdata[91 * 11 +  9] = 6'b001000;
assign fontdata[91 * 11 + 10] = 6'b000110;
assign fontdata[92 * 11 +  0] = 6'b000000;
assign fontdata[92 * 11 +  1] = 6'b001000;
assign fontdata[92 * 11 +  2] = 6'b001000;
assign fontdata[92 * 11 +  3] = 6'b001000;
assign fontdata[92 * 11 +  4] = 6'b001000;
assign fontdata[92 * 11 +  5] = 6'b001000;
assign fontdata[92 * 11 +  6] = 6'b001000;
assign fontdata[92 * 11 +  7] = 6'b001000;
assign fontdata[92 * 11 +  8] = 6'b001000;
assign fontdata[92 * 11 +  9] = 6'b001000;
assign fontdata[92 * 11 + 10] = 6'b000000;
assign fontdata[93 * 11 +  0] = 6'b110000;
assign fontdata[93 * 11 +  1] = 6'b001000;
assign fontdata[93 * 11 +  2] = 6'b001000;
assign fontdata[93 * 11 +  3] = 6'b001000;
assign fontdata[93 * 11 +  4] = 6'b001000;
assign fontdata[93 * 11 +  5] = 6'b000110;
assign fontdata[93 * 11 +  6] = 6'b001000;
assign fontdata[93 * 11 +  7] = 6'b001000;
assign fontdata[93 * 11 +  8] = 6'b001000;
assign fontdata[93 * 11 +  9] = 6'b001000;
assign fontdata[93 * 11 + 10] = 6'b110000;
assign fontdata[94 * 11 +  0] = 6'b000000;
assign fontdata[94 * 11 +  1] = 6'b000000;
assign fontdata[94 * 11 +  2] = 6'b000000;
assign fontdata[94 * 11 +  3] = 6'b000000;
assign fontdata[94 * 11 +  4] = 6'b010000;
assign fontdata[94 * 11 +  5] = 6'b101010;
assign fontdata[94 * 11 +  6] = 6'b000100;
assign fontdata[94 * 11 +  7] = 6'b000000;
assign fontdata[94 * 11 +  8] = 6'b000000;
assign fontdata[94 * 11 +  9] = 6'b000000;
assign fontdata[94 * 11 + 10] = 6'b000000;
assign fontdata[95 * 11 +  0] = 6'b000000;
assign fontdata[95 * 11 +  1] = 6'b000000;
assign fontdata[95 * 11 +  2] = 6'b000000;
assign fontdata[95 * 11 +  3] = 6'b011000;
assign fontdata[95 * 11 +  4] = 6'b111100;
assign fontdata[95 * 11 +  5] = 6'b111100;
assign fontdata[95 * 11 +  6] = 6'b011000;
assign fontdata[95 * 11 +  7] = 6'b000000;
assign fontdata[95 * 11 +  8] = 6'b000000;
assign fontdata[95 * 11 +  9] = 6'b000000;
assign fontdata[95 * 11 + 10] = 6'b000000;

endmodule
